module ROM_cost(
		d1_cntr,

		dw_1
	);

	localparam D1_IN_SIZE = 1;
	localparam D1_BW_W = 2;
	localparam D1_SHIFT = 0;
	localparam LOG2_D1_CYC = 9;
	localparam D1_CYC = 512;
	localparam D1_CH = 512;

	input [LOG2_D1_CYC-1:0] d1_cntr;

	output [D1_IN_SIZE*D1_BW_W-1:0] dw_1;

	reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_0 = { 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1 };

	assign dw_1 = dw_1_0[d1_cntr];

endmodule
